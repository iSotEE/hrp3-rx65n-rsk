/*
 *  TOPPERS/HRP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      High Reliable system Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tSIOPortCT11MPCore.cdl 285 2018-03-21 02:55:49Z ertl-hiro $
 */

/*
 *		シリアルインタフェースドライバのターゲット依存部（CT11MPCore用）
 *		のコンポーネント記述
 */

/*
 *  CT11MPcore with RealView Emulation Baseboard に関する定義
 */
import_C("ct11mpcore.h");

/*
 *  ARM PrimCell UART（PL011）用 簡易SIOドライバ
 */
import("tUartPL011.cdl");

/*
 *  シリアルインタフェースドライバのターゲット依存部の本体（シリアルイ
 *  ンタフェースドライバとSIOドライバを接続する部分）のセルタイプ
 */
celltype tSIOPortCT11MPCoreMain {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	[inline] entry		sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  SIOドライバとの結合
	 */
	call			sSIOPort	cSIOPort;
	[inline] entry	siSIOCBR	eiSIOCBR;

	/*
	 *  割込み要求ライン操作のための結合
	 */
	call	sInterruptRequest	cInterruptRequest;
};

/*
 *  シリアルインタフェースドライバのターゲット依存部（複合コンポーネン
 *  ト）のセルタイプ
 */
[active]
composite tSIOPortCT11MPCore {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	entry				sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  属性の定義
	 */
	attr {
		uintptr_t	baseAddress;				/* ベースアドレス */
		INTNO		interruptNumber;			/* 割込み番号 */
		PRI			isrPriority = 1;			/* ISR優先度 */
		PRI			interruptPriority = -2;		/* 割込み優先度 */

		uint8_t		ibrd = C_EXP("EB_UART_IBRD_38400");
		uint8_t		fbrd = C_EXP("EB_UART_FBRD_38400");
		uint8_t		lcr_h = C_EXP("UART_LCR_H_WLEN8");
	};

	/*
	 *  SIOドライバ
	 */
	cell tUartPL011 PL011 {
		baseAddress = composite.baseAddress;
		ibrd        = composite.ibrd;
		fbrd        = composite.fbrd;
		lcr_h       = composite.lcr_h;
		ciSIOCBR    = SIOPortMain.eiSIOCBR;
	};

	/*
	 *  シリアルインタフェースドライバのターゲット依存部の本体
	 */
	cell tSIOPortCT11MPCoreMain SIOPortMain {
		ciSIOCBR          => composite.ciSIOCBR;
		cSIOPort          = PL011.eSIOPort;
		cInterruptRequest = InterruptRequest.eInterruptRequest;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;

	/*
	 *  SIOの割込みサービスルーチンと割込み要求ライン
	 */
	cell tISR ISRInstance {
		interruptNumber = composite.interruptNumber;
		isrPriority     = composite.isrPriority;
		ciISRBody       = PL011.eiISR;
	};
	cell tInterruptRequest InterruptRequest {
		interruptNumber   = composite.interruptNumber;
		interruptPriority = composite.interruptPriority;
	};
};

/*
 *  これ以降のセルは，カーネルドメイン内に含める
 */
region rKernelDomain {

/*
 *  シリアルインタフェースドライバのターゲット依存部のプロトタイプ
 */
[prototype]
cell tSIOPortCT11MPCore SIOPortTarget1 {
	/* 属性の設定 */
	baseAddress     = C_EXP("EB_UART0_BASE");
	interruptNumber = C_EXP("EB_IRQNO_UART0");
};

[prototype]
cell tSIOPortCT11MPCore SIOPortTarget2 {
	/* 属性の設定 */
	baseAddress     = C_EXP("EB_UART1_BASE");
	interruptNumber = C_EXP("EB_IRQNO_UART1");
};

[prototype]
cell tSIOPortCT11MPCore SIOPortTarget3 {
	/* 属性の設定 */
	baseAddress     = C_EXP("EB_UART2_BASE");
	interruptNumber = C_EXP("EB_IRQN2_UART0");
};

[prototype]
cell tSIOPortCT11MPCore SIOPortTarget4 {
	/* 属性の設定 */
	baseAddress     = C_EXP("EB_UART3_BASE");
	interruptNumber = C_EXP("EB_IRQNO_UART3");
};
};
